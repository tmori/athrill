/*
 *		C言語で記述されたアプリケーションから，TECSベースのシリアルイン
 *		タフェースドライバを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id: tSerialAdapter.cdl 509 2016-01-12 06:06:14Z ertl-hiro $
 */
[singleton, active]
celltype tSerialAdapter {
	call	sSerialPort		cSerialPort[];
};
