/*
 *		C言語で記述されたアプリケーションから，TECSベースのテストプログ
 *		ラム用サービスを呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id: tTestServiceAdapter.cdl 884 2018-02-02 02:08:44Z ertl-hiro $
 */
[singleton, active]
celltype tTestServiceAdapter {
	call	sTestService	cTestService;
};
